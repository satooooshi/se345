module regfile( input logic clk, 
                input logic we3, 
                input logic [4:0] ra1, ra2, wa3, 
                input logic [31:0] wd3, 
                output logic [31:0] rd1, rd2);

    // logic [# of bits/word] rf[# of words(indicating address)]
    //Ex.
    //0x0:0x00000000
    //0x8:0x00000001
    //0x10:0x00000002
    logic [31:0] rf[31:0];

    //writeはwe3がHIの時のみ
    always_ff@(posedge clk)
        if(we3)rf[wa3]<=wd3;//rf[0x10]<=0x00000002

    //readはいつでも読み込まれる
    assign rd1=(ra1!=0)?rf[ra1]:0;
    assign rd2=(ra2!=0)?rf[ra2]:0;

endmodule