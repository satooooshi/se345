library verilog;
use verilog.vl_types.all;
entity calcutator_vlg_vec_tst is
end calcutator_vlg_vec_tst;
